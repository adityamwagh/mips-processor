module fullAdder_Dataflow(Cout, sum, in1, in2, Cin);
	input in1, in2;
	input Cin;
	output Cout;
	
	